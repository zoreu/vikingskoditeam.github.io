<?xml version="1.0" encoding="UTF-8" standalone="yes"?>

<channels>
	<!-- opicional -->
    <channels_info> <!-- this is opitonal -->
      <title>Para Amantes de Cinema</title> <!-- if channels_info, a title is required, other elements are optional -->
      <genre>News</genre>
      <description>this is the descripton string</description>
      <thumbnail>http://community-links.googlecode.com/svn/icons/news-icon.png</thumbnail>
      <fanart>http://community-links.googlecode.com/svn/icons/news-fanart.jpg</fanart>
      <date>20.10.2023</date>
      <credits>Gael</credits>
    </channels_info>
	<!-- opicional -->
    
    <channel>
        <name>Novo No Cine Room</name>
        <thumbnail>http://community-links.googlecode.com/svn/icons/news-icon.png</thumbnail>
        <fanart>http://community-links.googlecode.com/svn/icons/news-fanart.jpg</fanart>
		<info>Conteudos Recem-lançados no mundo</info>
		<externallink>http://localhost/gujal/itensrc.xml</externallink>
    </channel>
	
	<channel>
        <name>Populares</name>
        <thumbnail>http://community-links.googlecode.com/svn/icons/news-icon.png</thumbnail>
        <fanart>http://community-links.googlecode.com/svn/icons/news-fanart.jpg</fanart>
		<info>Filmes e series Populares</info>
		<externallink>https://bit.ly/3xZ2T9O</externallink>
    </channel>
	
   <channel>
        <name>Top Streaming</name>
        <thumbnail>http://community-links.googlecode.com/svn/icons/news-icon.png</thumbnail>
        <fanart>http://community-links.googlecode.com/svn/icons/news-fanart.jpg</fanart>
		<info>Filmes e Séries mais vistos em cada streaming</info>
		<externallink>https://bit.ly/3xZ2T9O</externallink>
   </channel>
   
   <channel>
        <name>Sagas</name>
        <thumbnail>http://community-links.googlecode.com/svn/icons/news-icon.png</thumbnail>
        <fanart>http://community-links.googlecode.com/svn/icons/news-fanart.jpg</fanart>
		<info>Melhores coletaneas</info>
		<externallink>https://bit.ly/3xZ2T9O</externallink>
   </channel>
   
   <channel>
        <name>Melhor Avaliação</name>
        <thumbnail>http://community-links.googlecode.com/svn/icons/news-icon.png</thumbnail>
        <fanart>http://community-links.googlecode.com/svn/icons/news-fanart.jpg</fanart>
		<info>Filmes e Séries mais bem avaliados</info>
		<externallink>https://bit.ly/3xZ2T9O</externallink>
   </channel>

</channels>	